library ieee;
use ieee.std_logic_1164.all;

entity REG is
    port (
        instrucao_in : in std_logic_vector(7 downto 0);
        instrucao_out : out std_logic_vector(2 downto 0)
    );
end entity REG;

architecture behavioral of REG is
begin

	 
end architecture behavioral;